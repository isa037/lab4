library ieee;
use ieee.numeric_std.all;
USE IEEE.STD_LOGIC_1164.ALL;


package my_pkg is
  type array33 is array (natural range <>) of std_logic_vector(32 downto 0);
  type array36 is array (natural range <>) of std_logic_vector(35 downto 0);
end package;

package body my_pkg is
end package body;
