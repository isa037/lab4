LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FFN_EN_FP IS
	PORT (R : IN STD_LOGIC;
			ENABLE, CLOCK, RESETN : IN STD_LOGIC;
			Q :	OUT STD_LOGIC);
END FFN_EN_FP;

ARCHITECTURE BEHAVIOR OF FFN_EN_FP IS
BEGIN
	PROCESS (CLOCK, RESETN)
	BEGIN
		IF (RESETN = '0') THEN   -- RST ASINCRONO ATTIVO BASSO
			Q <= '0';
		ELSIF (CLOCK'EVENT AND CLOCK = '1') THEN
			IF ENABLE='1' THEN
				Q <= R;
			END IF;
		END IF;
	END PROCESS;
END BEHAVIOR;
